module MAS16bA (
        input clk
);

endmodule
